module fifo #(

) (

);

endmodule
